/*
 * @Author      : myyerrol
 * @Date        : 2024-11-02 15:22:27
 * @LastEditors : myyerrol
 * @LastEditTime: 2024-11-02 15:24:04
 * @Description : First Input First Out
 *
 * Copyright (c) 2024 by MEMDSL, All Rights Reserved.
 */

module fifo #(
    parameter DATA_WIDTH = 32
) (
    input logic i_clk,
    input logic i_rst_n,

);

endmodule
