/*
 * @Author      : myyerrol
 * @Date        : 2024-11-01 20:01:17
 * @LastEditors : myyerrol
 * @LastEditTime: 2024-12-26 11:01:34
 * @Description : Register defines.
 *
 * Copyright (c) 2024 by MEMDSL, All Rights Reserved.
 */

`define REG_DELAY_CYCLE 0
