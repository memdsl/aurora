/*
 * @Author      : myyerrol
 * @Date        : 2024-11-01 20:01:17
 * @LastEditors : myyerrol
 * @LastEditTime: 2024-11-02 15:20:06
 * @Description : Configs.
 *
 * Copyright (c) 2024 by MEMDSL, All Rights Reserved.
 */

`define DELAY_CYCLE 0
