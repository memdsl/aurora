`define DELAY_CYCLE 0
