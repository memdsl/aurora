/*
 * @Author      : myyerrol
 * @Date        : 2024-07-02 12:49:46
 * @LastEditors : myyerrol
 * @LastEditTime: 2024-07-07 22:30:11
 * @FilePath    : /memdsl/aurora/src/sv/common/mul/rtl/mul_nnbit_shift.sv
 * @Description : nnbit shift multiplier
 *
 * Copyright (c) 2024 by myyerrol, All Rights Reserved.
 */

module mul_nnbit_shift #(
    parameter DATA_WIDTH = 8
) (
    input  logic                          i_clk,
    input  logic                          i_rst_n,
    input  logic [DATA_WIDTH - 1     : 0] i_num_x,
    input  logic [DATA_WIDTH - 1     : 0] i_num_y,
    output logic                          o_end,
    output logic [DATA_WIDTH * 2 - 1 : 0] o_res
);

    logic [DATA_WIDTH * 2 - 1 : 0] r_num_x;
    logic [DATA_WIDTH     - 1 : 0] r_num_y;
    logic [DATA_WIDTH * 2 - 1 : 0] r_res;

    logic [DATA_WIDTH * 2 - 1 : 0] w_res;

    int count;

    always_ff @(posedge i_clk) begin
        if (!i_rst_n) begin
            r_num_x <= {{DATA_WIDTH{i_num_x[DATA_WIDTH - 1]}}, i_num_x};
            r_num_y <= i_num_y;
            r_res   <= {(DATA_WIDTH * 2){1'b0}};
            count   <= 0;
        end
        else begin
            if (count == DATA_WIDTH) begin
                o_end <= 1'b1;
                o_res <= r_res + (~w_res + 1'b1);
                count <= count;
            end
            else begin
                o_end   <= 1'b0;
                o_res   <= {(DATA_WIDTH * 2){1'b0}};
                r_res   <= r_res + w_res;
                r_num_x <= (r_num_x << 1);
                r_num_y <= (r_num_y >> 1);
                count   <= count + 1'b1;
            end
        end
    end

    assign w_res = (r_num_y[0]) ? r_num_x : {(DATA_WIDTH * 2){1'b0}};

endmodule
